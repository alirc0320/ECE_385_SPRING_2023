//module background_collision_example (
//	input logic [9:0] DrawX, DrawY,
//	input logic vga_clk, blank,
//	output logic [3:0] red, green, blue
//);
//
//logic [17:0] rom_address;
//logic [3:0] rom_q;
//
//logic [3:0] palette_red, palette_green, palette_blue;
//
//assign rom_address = ((DrawX * 500) / 640) + (((DrawY * 500) / 480) * 500);
//
//always_ff @ (posedge vga_clk) begin
//	red <= 4'h0;
//	green <= 4'h0;
//	blue <= 4'h0;
//
//	if (blank) begin
//		red <= palette_red;
//		green <= palette_green;
//		blue <= palette_blue;
//	end
//end
//
//background_collision_rom background_collision_rom (
//	.clock   (vga_clk),
//	.address (rom_address),
//	.q       (rom_q)
//);
//
//background_collision_palette background_collision_palette (
//	.index (rom_q),
//	.red   (palette_red),
//	.green (palette_green),
//	.blue  (palette_blue)
//);
//
//endmodule
